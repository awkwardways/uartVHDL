library ieee;
use ieee.std_logic_1164.all;

entity tx is 
  port(
    txLine        : out std_logic := '1';
    parallelIn    : in std_logic_vector(7 downto 0);
    loadTransmit  : in std_logic;
    baudIn        : in std_logic
  );
end entity tx;

architecture rtl of tx is 
  type transmissionState is (idle, startBit, stopBit, data);
  signal currentState : transmissionState := idle;
  signal byteBuffer   : std_logic_vector(7 downto 0) := x"00";

begin

  loadByte: process(baudIn)
  begin
    if rising_edge(baudIn) then
      if loadTransmit = '1' then
        byteBuffer <= parallelIn;
      end if;
    end if;
  end process loadByte;  

  transmitByte: process(baudIn)
    variable isTransmitting : std_logic := '0';
    variable currentBit : natural := 0; 
    -- variable coolDown : integer := 0;
  begin
    if rising_edge(baudIn) then

      if loadTransmit = '0' then -- if loadTransmit = '0' and coolDown >= 9599 then
        isTransmitting := '1';
        -- coolDown := 0;
      -- else
        -- isTransmitting := '0';
        -- coolDown := coolDown + 1;
      end if;

      case currentState is
        when idle =>
          txLine <= not isTransmitting;
          currentState <= startBit;
          if isTransmitting = '0' then
            currentState <= idle;
          end if;
        
        when startBit =>
          currentState <= data;
          txLine <= byteBuffer(currentBit);
          currentBit := currentBit + 1;
        
        when data =>
          if currentBit = 8 then
            txLine <= '1';
            currentBit := 0;
            currentState <= stopBit;
          else
            txLine <= byteBuffer(currentBit);
            currentBit := currentBit + 1;
          end if;
            
        
        when stopBit =>
          currentState <= idle;
          isTransmitting := '0';
      end case;
    end if;
  end process;

end architecture;